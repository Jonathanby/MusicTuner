`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:13:38 11/08/2016 
// Design Name: 
// Module Name:    Cap_Note 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Cap_Note(
    );


/*
	all new shiz
	should i use the built in a to d converter
	or will the signal from the key would be enough
	test latter first with gen_note, then actual note
*/

endmodule
