`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:49:42 11/08/2016 
// Design Name: 
// Module Name:    Listen_Graph 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Listen_Graph(
    );
	 
	 //input x and y
	 //output rgb hsync vsync?

//for listen button and listen box
//listen mode box
//and listen frequency box

//hilight or not hilight mode


endmodule
